//Verilog HDL for "Lab3", "Inverter" "functional"

`timescale 1ns/10ps

module Inverter ( Vout, Vin );

  input Vin;
  output Vout;

  not #1 n1(Vout,Vin);	

endmodule
